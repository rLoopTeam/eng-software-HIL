`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:02:31 03/26/2016 
// Design Name: 
// Module Name:    SimplePodModel 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module SimplePodModel(
    input [31:0] accel,
    input clk_200khz,
    output [31:0] position,
    output [31:0] velocity
    );


endmodule
